module ps2_decoder(
    input wire clk,

    input wire ps2_clk,
    input wire ps2_data,

    output logic [7:0] data
    );

    // your code goes here!
    assign data = 0;

endmodule